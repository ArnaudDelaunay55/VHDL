LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

PACKAGE ONDES_PKG IS
TYPE TABLEAU IS ARRAY (NATURAL RANGE <>) OF NATURAL;
CONSTANT SINUS_ROM : TABLEAU :=(
0	,
6	,
13	,
19	,
25	,
31	,
38	,
44	,
50	,
56	,
63	,
69	,
75	,
81	,
88	,
94	,
100	,
106	,
112	,
118	,
124	,
130	,
137	,
143	,
149	,
155	,
161	,
167	,
172	,
178	,
184	,
190	,
196	,
202	,
207	,
213	,
219	,
225	,
230	,
236	,
241	,
247	,
252	,
258	,
263	,
269	,
274	,
279	,
284	,
290	,
295	,
300	,
305	,
310	,
315	,
320	,
325	,
330	,
334	,
339	,
344	,
348	,
353	,
358	,
362	,
366	,
371	,
375	,
379	,
384	,
388	,
392	,
396	,
400	,
404	,
407	,
411	,
415	,
419	,
422	,
426	,
429	,
433	,
436	,
439	,
442	,
445	,
449	,
452	,
454	,
457	,
460	,
463	,
465	,
468	,
471	,
473	,
475	,
478	,
480	,
482	,
484	,
486	,
488	,
490	,
492	,
493	,
495	,
497	,
498	,
500	,
501	,
502	,
503	,
504	,
505	,
506	,
507	,
508	,
509	,
510	,
510	,
511	,
511	,
511	,
512	,
512	,
512	

);
END PACKAGE ONDES_PKG;
